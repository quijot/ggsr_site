Nombre:      david gonzalez
Correo:      david.gonzalez@anda.gob.sv
Institucion: anda
Direccion:   san miguel
Ciudad/Pais: san miguel, el salvador 
Telefono:    2600 2600
Descripcion: 
